* C:\Users\User\Desktop\lab simulate file\lab 7.sch

* Schematics Version 9.1 - Web Update 1
* Sat Sep 26 23:34:43 2020


.PARAM         RVAR=10 

** Analysis setup **
.DC LIN PARAM RVAR 1 20 0.1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "lab 7.net"
.INC "lab 7.als"


.probe


.END
